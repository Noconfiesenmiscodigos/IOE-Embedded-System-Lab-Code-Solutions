--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   11:48:23 02/26/2022
-- Design Name:   
-- Module Name:   D:/Lab_2/Multiplexer/Demultiplexer_TB.vhd
-- Project Name:  Multiplexer
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Demultiplexer
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY Demultiplexer_TB IS
END Demultiplexer_TB;
 
ARCHITECTURE behavior OF Demultiplexer_TB IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Demultiplexer
    PORT(
         A : IN  std_logic;
         S : IN  std_logic_vector(1 downto 0);
         Y : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal A : std_logic := '0';
   signal S : std_logic_vector(1 downto 0) := (others => '0');

 	--Outputs
   signal Y : std_logic_vector(3 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant <clock>_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Demultiplexer PORT MAP (
          A => A,
          S => S,
          Y => Y
        );

   -- Clock process definitions
  -- <clock>_process :process
   --begin
		--<clock> <= '0';
		--wait for <clock>_period/2;
		--<clock> <= '1';
		--wait for <clock>_period/2;
   --end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

     -- wait for <clock>_period*10;

      -- insert stimulus here 
		
		A<='1';
		S<="00";
		wait for 100 ns;
		S<="01";
		wait for 100 ns;
		S<="10";
		wait for 100 ns;
		S<="11";
		
		A<='0';
		S<="00";
		wait for 100 ns;
		S<="01";
		wait for 100 ns;
		S<="10";
		wait for 100 ns;
		S<="11";

      wait;
   end process;

END;
